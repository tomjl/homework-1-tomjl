module sum_prod_tb;

  // complete the testbench

endmodule;

module multiplier (
  input  logic [15:0]a,b,
  output logic [31:0] product
);

// complete the module

endmodule

module sum_prod #(parameter N) (
  input  logic [N-1:0] X [5:0],
  output logic [2N+2:0] result
);

// complete the module

endmodule

module multiplier #(parameter N) (
  input  logic [N-1:0]a,b,
  output logic [2*N-1:0] product
);

// complete the module

endmodule

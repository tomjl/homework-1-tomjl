module multiplier_tb;

  // complete

endmodule

module multiplier_tb;

  localparam N = 4;

  // complete
endmodule

module count_1 (
  input logic [3:0] a,
  output logic [2:0] out
);
  // …
  // Add your description here
  // …
endmodule

module bin2gray (
  input logic [3:0] binary,
  output logic [3:0] gray
);
  // …
  // Add your description here
  // …
endmodule
